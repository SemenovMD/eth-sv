package pkg_tb;


    
endpackage